`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   14:36:39 09/16/2016
// Design Name:   ALU_Decoder
// Module Name:   C:/xilingProjects/Lab3_ControlUnit/ALU_Decoder_TestFixture.v
// Project Name:  Lab3_ControlUnit
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: ALU_Decoder
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module ALU_Decoder_TestFixture;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	ALU_Decoder uut (
		.()
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

