`timescale 1ns / 1ps

module ControlUnit_VerilogModule(  ALU_Decoder);


endmodule
